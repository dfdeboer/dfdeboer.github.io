A circuit with two op-amps
*
***************MAIN CIRCUIT************
*      From  To    From  To     <--(for current sources)
*Part  or    or    or    or
*Name  +     -     +     -     value
R1     2     0                 20kohms
R2     2     4                 20kohms
R3     1     3                 15kohms
R4     5     3                 30kohms
R5     4     5                 50khoms
X1     2     1     4           uA741_op_amp
X2     3     0     5           uA741_op_amp
VS     1     0                 2.5volts
*
***************SUB CIRCUIT************
*The op-amp model follows:
.subckt uA741_op_amp                  1  2  4
* Connections:                        |  |  |
*     Node 1 is the inverting input---+  |  |
*     Node 2 is the non-inverting input--+  |
*     Node 4 is the output------------------+
*
Gm     0     3     2     1     0.2msiemens
R1     3     0                 1Gohm
C1     3     0                 30pf
Eout   4     0     3     0     1
Iopen1 0     1                 0amps
Iopen2 0     2                 0amps
.ends uA741_op_amp
*
.end

