An op-amp circuit with a model of a uA741 op-amp included
*
***************MAIN CIRCUIT************
*      From  To    From  To     <--(for current sources)
*Part  or    or    or    or
*Name  +     -     +     -     value
Rf     4     1                 10kohms
Rin    5     1                 1kohm
X1     1     2     4           uA741_op_amp
*                 (^connect op-amp output to node 4)
* Elements added to provide stimulus and response
Vin    5     0                 1volt
V0     2     0                 0volts
Rload  4     0                 1kohm
*
***************SUB CIRCUIT************
*The op-amp model follows:
.subckt uA741_op_amp                  1  2  4
* Connections:                        |  |  |
*     Node 1 is the inverting input---+  |  |
*     Node 2 is the non-inverting input--+  |
*     Node 4 is the output------------------+
*
Gm     0     3     2     1     0.2msiemens
R1     3     0                 1Gohm
C1     3     0                 30pf
Eout   4     0     3     0     1
Iopen1 0     1                 0amps
Iopen2 0     2                 0amps
.ends uA741_op_amp
*
.end

