*-------------------------------------------------------------------------------
*                    TN0606 n-ch Enhancement MOSFET (model from Supertex)
.MODEL TN0606   NMOS (LEVEL=3       RS=0.100        NSUB=3.00E15    DELTA=0.1
+                    KAPPA=0.10123  TPG=1           CGDO=4.3432E-11 RD=0.45
+                    VTO=1.300      VMAX=1.0E7      ETA=0.0223089   NFS=6.6E10
+                    TOX=1.00E-7    LD=1.698E-9     UO=862.425      XJ=6.46E-7
+                    THETA=1.0E-5   CGSO=1.2179E-10 L=2.5E-6        W=2.0E-2)
*-------------------------------------------------------------------------------
*                    TP0606 p-ch Enhancement MOSFET (model from Supertex)
.MODEL TP0606   PMOS (LEVEL=3       RS=0.200        NSUB=3.00E15    DELTA=0.1
+                    KAPPA=0.0821   TPG=-1          CGDO=5.2212E-11 RD=0.854
+                    VTO=-2.100     VMAX=3.0E6      ETA=0.12098     NFS=3.384E11
+                    TOX=1.00E-7    LD=1.1400E-9    UO=365.45       XJ=6.5E-7
+                    THETA=4.063E-5 CGSO=8.532E-11  L=2.5E-6        W=2.0E-2)

